-- Ocupo que este componente haga lo siguiente
    -- Estados que manejen la secuencia de pasos