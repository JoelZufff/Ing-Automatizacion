process(entrada_num)
	begin
		case