library	IEEE;
use	IEEE.std_logic_1164.all;	 

entity Maquina_expendedora is
    port 
    (
        CLK     : in std_logic;
        RST     : in std_logic;
           
    );
end entity;

architecture Venta of Maquina_expendedora is
begin

    -- Establecer el reloj de cambio de estado
    -- 

end Venta;